//Main will connect the keyboard to the actual program
module main();
endmodule
