module pearson_hash8(message, reset_n, random_table, hash, counter);
	//Assume 8 bit wide sequencing
	input [7:0] message;
	input reset_n;
	output [7:0] hash;
	output reg [2:0] counter = 3'b000;
	
	//Intialize variables for computation
	reg [7:0] temp_hash = 7'b0;
	reg [7:0] access_point;
	
	//Loop over 8 bits of input
	always @(*) begin
		if (!reset_n)
			temp_hash <= 7'b0;
			access_point <= 7'b0;
			counter <= 3'b000;
			
		else if (counter != 3'b111) begin
			access_point <= temp_hash ^ message; 
			temp_hash <= random_table[access_point: (access_point + 8)];
			counter <= counter + 1;
		end
	end
	
	//Output final sequenceof bits
	assign hash = (counter == 3'b111) ? temp_hash : 8'b0;
endmodule