`include "../Hash/pearson_hash8.v"

module make_starting_memory(starting_memory);
	output [47:0] starting_memory;
	
	wire p1_money = 8'b00110010;
	wire p2_money = 8'b00110010;
	wire p1_private = 8'b01110101;
	wire p2_private = 8'b00011011;
	
endmodule