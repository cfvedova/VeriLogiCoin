module store_values()
	if(process == 3'b100)
endmodule